// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	LandminesBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input	logic	SingleHitPulse,

					output	logic	drawingRequest_mine1, //output that the pixel should be dispalyed
					output	logic	drawingRequest_mine2, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 

logic mine1_flag;
logic mine2_flag;

logic [0:14] [0:16] [3:0] MazeBitMapMask = 
{	
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00}
};


logic [0:1] [0:31] [0:31] [7:0]  object_colors  = {
	// LANDMINE - MINE TYPE 1 ( 01 CODE )
   {{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h91,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hb6,8'h6d,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'h6d,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hb6,8'h24,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hb6,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hda,8'h8d,8'h60,8'h80,8'ha4,8'hc4,8'hcd,8'hb1,8'hb6,8'hb6,8'hb6,8'h6d,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb1,8'hf1,8'hc0,8'hc0,8'hc0,8'hc0,8'ha0,8'h80,8'h64,8'h91,8'hd6,8'h91,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hcd,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'ha0,8'h84,8'h91,8'hda,8'h91,8'h24,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf1,8'hc0,8'he0,8'he0,8'he0,8'he0,8'hc0,8'hc0,8'ha0,8'had,8'hd6,8'hb6,8'h6d,8'h24,8'h6d,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hb6,8'hd1,8'hc0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hc0,8'hc0,8'hc4,8'hb1,8'h6d,8'h24,8'h24,8'h6d,8'hb1,8'h8d,8'hb6,8'hda,8'hda,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'h91,8'h6d,8'h8d,8'hc0,8'he0,8'he0,8'he0,8'he4,8'he4,8'he4,8'he4,8'he0,8'hc0,8'hc0,8'ha4,8'h64,8'h24,8'h24,8'h6d,8'h8d,8'h60,8'h24,8'h24,8'h24,8'hb6,8'hff,8'hff},
	{8'hff,8'hff,8'hb6,8'hb6,8'hda,8'hff,8'hff,8'hd1,8'hc0,8'he0,8'he0,8'he4,8'hed,8'hed,8'hed,8'he4,8'he4,8'hc0,8'hc0,8'ha0,8'h80,8'h80,8'h60,8'h64,8'h80,8'h80,8'h60,8'h24,8'h91,8'hda,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hb6,8'h6d,8'h91,8'hda,8'hcd,8'he0,8'he0,8'he4,8'he4,8'hed,8'hed,8'hed,8'he5,8'he4,8'hc0,8'ha0,8'ha0,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h84,8'h8d,8'hb6,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hb6,8'h24,8'h64,8'hc0,8'hc0,8'he0,8'he4,8'he4,8'hed,8'hed,8'hed,8'hed,8'he4,8'hc0,8'h84,8'h64,8'h24,8'h60,8'h60,8'h80,8'h60,8'h80,8'ha4,8'hb1,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h84,8'hc0,8'hc0,8'he0,8'he4,8'he4,8'hed,8'hed,8'hed,8'he4,8'hc4,8'h84,8'h6d,8'h25,8'h24,8'h24,8'h20,8'h60,8'h60,8'h80,8'had,8'hd1,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hcd,8'hc0,8'hc0,8'he0,8'he0,8'he4,8'he4,8'he4,8'he4,8'he4,8'ha4,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h64,8'h60,8'h60,8'had,8'hd1,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hd1,8'hc0,8'hc0,8'hc0,8'he0,8'he0,8'he4,8'he4,8'he4,8'hc0,8'h84,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h64,8'h60,8'h60,8'ha4,8'hd1,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'had,8'ha0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h64,8'h60,8'h60,8'ha4,8'had,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h91,8'hb1,8'ha0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'ha0,8'ha0,8'h80,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h60,8'h60,8'h60,8'h80,8'h84,8'hb6,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hb6,8'h92,8'hb6,8'ha5,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'h60,8'h24,8'h24,8'h65,8'h8d,8'h64,8'h60,8'h60,8'h80,8'h80,8'h24,8'h24,8'hb6,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hb6,8'h91,8'h91,8'h6d,8'h64,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'h80,8'h80,8'h80,8'h60,8'h84,8'h84,8'h80,8'h80,8'h80,8'h80,8'had,8'h91,8'h91,8'h91,8'hda,8'hff},
	{8'hff,8'hff,8'hda,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h80,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'h80,8'h80,8'h80,8'h80,8'h80,8'ha0,8'ha0,8'ha0,8'h80,8'h80,8'ha4,8'hd6,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h80,8'h80,8'h80,8'h80,8'had,8'hd6,8'had,8'h80,8'h80,8'ha0,8'ha4,8'ha4,8'hc4,8'ha4,8'ha0,8'ha0,8'hd1,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hd6,8'ha4,8'h80,8'h64,8'hb6,8'hff,8'hb6,8'h24,8'h20,8'h84,8'hc4,8'hcd,8'hed,8'hc5,8'hc4,8'hd1,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hd6,8'had,8'h64,8'h91,8'hff,8'h91,8'h24,8'h00,8'h64,8'hcd,8'hed,8'hed,8'ha4,8'hb1,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h91,8'h91,8'hff,8'h91,8'h24,8'h20,8'h84,8'ha4,8'had,8'hb1,8'h6d,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h91,8'hda,8'h6d,8'h24,8'h65,8'hb1,8'h8d,8'h6d,8'hb2,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h91,8'hd6,8'h24,8'h24,8'hb6,8'hff,8'hff,8'h91,8'h91,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'h24,8'h91,8'hff,8'hff,8'hff,8'hff,8'hda,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h91,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h91,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}}
	,// TNT - MINE TYPE 2 ( 02 CODE )
   {{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hcd,8'had,8'had,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb1,8'hb1,8'hff,8'hff,8'hff,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hcd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf1,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb1,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hec,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hed,8'he4,8'hff,8'hff,8'hff,8'hb1,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hff,8'hff,8'hec,8'hff,8'hff,8'hec,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hf6,8'hed,8'hed,8'he4,8'hf1,8'hed,8'hed,8'hc5,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hd1,8'hff,8'hed,8'hec,8'hec,8'hec,8'hf1,8'hec,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hf5,8'hed,8'hed,8'he4,8'hf1,8'hed,8'hed,8'he4,8'hfa,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hec,8'hec,8'hf8,8'hf8,8'hec,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hed,8'hed,8'hed,8'he4,8'hed,8'hed,8'hed,8'he4,8'hed,8'hed,8'hed,8'hff,8'hff,8'hff,8'hff,8'hff,8'hec,8'hec,8'hec,8'hec,8'hf8,8'hf8,8'hf8,8'hec,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h6d,8'h96,8'h6d,8'h6d,8'h6d,8'h6d,8'had,8'hed,8'hed,8'hed,8'hed,8'hed,8'hcc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hec,8'hec,8'hf8,8'hec,8'hf4,8'hec,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h6d,8'hb6,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hed,8'hed,8'he4,8'hcd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hec,8'hff,8'hec,8'hff,8'hf6,8'hec,8'hec,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hf6,8'hed,8'hed,8'h85,8'hfe,8'hfd,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hec,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hed,8'hed,8'hec,8'hfd,8'hf8,8'hfc,8'hfc,8'hfd,8'h6d,8'h24,8'h24,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hed,8'hed,8'hec,8'hfd,8'hfc,8'h6d,8'hf8,8'hfc,8'hf8,8'he5,8'h25,8'h24,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hf5,8'hed,8'hfd,8'hfc,8'hfc,8'hd4,8'hb5,8'hfd,8'hfc,8'hf8,8'hed,8'hc4,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hf5,8'hed,8'hfd,8'hfc,8'hf8,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hed,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hed,8'hed,8'hfc,8'hfc,8'hf8,8'hfc,8'h6d,8'hf8,8'hfc,8'hfc,8'hed,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hed,8'hed,8'hed,8'hfc,8'hfc,8'hfd,8'h6d,8'hfd,8'hfc,8'hfc,8'hf8,8'hed,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hf6,8'hed,8'hed,8'hfc,8'hf8,8'h64,8'hfc,8'hfc,8'hfc,8'hfc,8'hc4,8'hc4,8'hf1,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'h6d,8'hed,8'hed,8'hf8,8'hfc,8'h6c,8'h6d,8'hfc,8'hfc,8'hf8,8'he4,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hb6,8'h91,8'h6d,8'hfd,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hc4,8'hed,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'he5,8'h96,8'h6d,8'h6d,8'h6d,8'hfc,8'hfc,8'hfc,8'hfc,8'hec,8'hed,8'hed,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hf5,8'hed,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6c,8'h6d,8'h24,8'h24,8'h24,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hf5,8'hed,8'hed,8'hc4,8'h6d,8'h6d,8'h91,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hed,8'hed,8'hed,8'he4,8'hf1,8'hed,8'hf1,8'h8d,8'h6d,8'h24,8'h24,8'h64,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hf6,8'hed,8'he4,8'hed,8'hed,8'hed,8'hed,8'he4,8'hed,8'hed,8'hed,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hf1,8'hed,8'hed,8'he4,8'hed,8'hed,8'hed,8'he4,8'hf6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hc4,8'hcd,8'hff,8'hed,8'hed,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}}
 };
			


// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask <= 
{	
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00}
};
	end
	else begin
	   // default values
		RGBout <= TRANSPARENT_ENCODING ;
		mine1_flag <= 1'b0;
		mine2_flag <= 1'b0;
		
	
		if (InsideRectangle == 1'b1 ) begin // take bits 5,6,7,8,9,10 from address to select  position in the maze
			
			// type 1 mine
		   if (MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h01)   
				begin
						RGBout <= object_colors[0][offsetY[4:0]][offsetX[4:0]] ;
						mine1_flag <= 1'b1;
				end
		
		// type 2 mine
			else if (MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h02)
				begin
						RGBout <= object_colors[1][offsetY[4:0]][offsetX[4:0]] ;
						mine2_flag <= 1'b1;
				end
				
			 if (SingleHitPulse)
					MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h00;
	
		end
	end
		
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest_mine1 = ( (RGBout != TRANSPARENT_ENCODING ) && mine1_flag ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmap
assign drawingRequest_mine2 = ( (RGBout != TRANSPARENT_ENCODING ) && mine2_flag ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmap   
endmodule

